xml.instruct! :xml, :version => "1.0"

xml.status do
  xml.result 'success'
end
